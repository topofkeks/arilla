-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Sat Aug 21 02:42:49 2021"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY SevenSegmentInterface1 IS 
	PORT
	(
		bit0 :  IN  STD_LOGIC;
		bit1 :  IN  STD_LOGIC;
		bit2 :  IN  STD_LOGIC;
		bit3 :  IN  STD_LOGIC;
		b :  OUT  STD_LOGIC;
		c :  OUT  STD_LOGIC;
		d :  OUT  STD_LOGIC;
		e :  OUT  STD_LOGIC;
		f :  OUT  STD_LOGIC;
		g :  OUT  STD_LOGIC;
		dp :  OUT  STD_LOGIC;
		a :  OUT  STD_LOGIC
	);
END SevenSegmentInterface1;

ARCHITECTURE bdf_type OF SevenSegmentInterface1 IS 

SIGNAL	NOTbit0 :  STD_LOGIC;
SIGNAL	NOTbit1 :  STD_LOGIC;
SIGNAL	NOTbit2 :  STD_LOGIC;
SIGNAL	NOTbit3 :  STD_LOGIC;
SIGNAL	one :  STD_LOGIC;
SIGNAL	zero :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;


BEGIN 



NOTbit0 <= NOT(bit0);



NOTbit1 <= NOT(bit1);



SYNTHESIZED_WIRE_3 <= NOTbit0 AND bit2;


SYNTHESIZED_WIRE_4 <= bit1 AND bit2;


SYNTHESIZED_WIRE_5 <= NOTbit1 AND NOTbit3;


SYNTHESIZED_WIRE_35 <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4 OR SYNTHESIZED_WIRE_5;


SYNTHESIZED_WIRE_6 <= NOTbit0 AND NOTbit2 AND NOTbit3;


SYNTHESIZED_WIRE_8 <= NOTbit0 AND bit2 AND bit3;


SYNTHESIZED_WIRE_7 <= bit0 AND NOTbit2 AND bit3;


SYNTHESIZED_WIRE_9 <= NOTbit1 AND NOTbit2;


SYNTHESIZED_WIRE_10 <= NOTbit1 AND NOTbit3;


SYNTHESIZED_WIRE_36 <= SYNTHESIZED_WIRE_6 OR SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10 OR zero;


NOTbit2 <= NOT(bit2);





SYNTHESIZED_WIRE_11 <= NOTbit0 AND NOTbit2;


SYNTHESIZED_WIRE_13 <= NOTbit0 AND bit3;


SYNTHESIZED_WIRE_12 <= NOTbit2 AND bit3;


SYNTHESIZED_WIRE_14 <= NOTbit0 AND bit1;


SYNTHESIZED_WIRE_15 <= bit0 AND NOTbit1;


SYNTHESIZED_WIRE_37 <= SYNTHESIZED_WIRE_11 OR SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15 OR zero;


SYNTHESIZED_WIRE_16 <= NOTbit0 AND NOTbit1 AND NOTbit3;


NOTbit3 <= NOT(bit3);



SYNTHESIZED_WIRE_18 <= NOTbit1 AND bit2 AND bit3;


SYNTHESIZED_WIRE_17 <= bit1 AND NOTbit2 AND bit3;


SYNTHESIZED_WIRE_19 <= bit1 AND bit2 AND NOTbit3;


SYNTHESIZED_WIRE_20 <= bit0 AND NOTbit2;


SYNTHESIZED_WIRE_38 <= SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17 OR SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20 OR zero;


SYNTHESIZED_WIRE_21 <= NOTbit1 AND NOTbit3;


SYNTHESIZED_WIRE_24 <= bit2 AND NOTbit3;


SYNTHESIZED_WIRE_22 <= bit0 AND bit2;


SYNTHESIZED_WIRE_23 <= bit0 AND bit1;


SYNTHESIZED_WIRE_39 <= SYNTHESIZED_WIRE_21 OR SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23 OR SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_25 <= NOTbit0 AND bit1 AND NOTbit2;


SYNTHESIZED_WIRE_27 <= NOTbit2 AND NOTbit3;


SYNTHESIZED_WIRE_26 <= bit1 AND NOTbit3;


SYNTHESIZED_WIRE_28 <= bit0 AND NOTbit1;


SYNTHESIZED_WIRE_29 <= bit0 AND bit2;


SYNTHESIZED_WIRE_40 <= SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27 OR SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29 OR zero;


SYNTHESIZED_WIRE_30 <= NOTbit0 AND bit1 AND NOTbit2;


SYNTHESIZED_WIRE_32 <= NOTbit1 AND bit2;


SYNTHESIZED_WIRE_31 <= bit2 AND NOTbit3;


SYNTHESIZED_WIRE_33 <= bit0 AND NOTbit1;


SYNTHESIZED_WIRE_34 <= bit0 AND bit3;


SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_31 OR SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_34 OR zero;


a <= NOT(SYNTHESIZED_WIRE_35);



b <= NOT(SYNTHESIZED_WIRE_36);



c <= NOT(SYNTHESIZED_WIRE_37);



d <= NOT(SYNTHESIZED_WIRE_38);



e <= NOT(SYNTHESIZED_WIRE_39);



f <= NOT(SYNTHESIZED_WIRE_40);



g <= NOT(SYNTHESIZED_WIRE_41);



SYNTHESIZED_WIRE_0 <= bit0 AND NOTbit1 AND NOTbit2;


SYNTHESIZED_WIRE_2 <= NOTbit0 AND bit1 AND bit3;


SYNTHESIZED_WIRE_1 <= bit0 AND NOTbit3;

dp <= one;

one <= '1';
zero <= '0';
END bdf_type;