-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Mon Aug 30 00:51:18 2021"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY SRAMAdapter IS 
	PORT
	(
		RD :  IN  STD_LOGIC;
		WR :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		ADDR :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		ByteEnable :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA :  INOUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END SRAMAdapter;

ARCHITECTURE bdf_type OF SRAMAdapter IS 

COMPONENT sram32_arilla
	PORT(wren : IN STD_LOGIC;
		 rden : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
		 byteena : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	HIT :  STD_LOGIC;
SIGNAL	rden :  STD_LOGIC;
SIGNAL	wren :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	DFF_inst3 :  STD_LOGIC;


BEGIN 



PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(31) <= SYNTHESIZED_WIRE_0(31);
ELSE
	DATA(31) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(30) <= SYNTHESIZED_WIRE_0(30);
ELSE
	DATA(30) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(29) <= SYNTHESIZED_WIRE_0(29);
ELSE
	DATA(29) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(28) <= SYNTHESIZED_WIRE_0(28);
ELSE
	DATA(28) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(27) <= SYNTHESIZED_WIRE_0(27);
ELSE
	DATA(27) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(26) <= SYNTHESIZED_WIRE_0(26);
ELSE
	DATA(26) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(25) <= SYNTHESIZED_WIRE_0(25);
ELSE
	DATA(25) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(24) <= SYNTHESIZED_WIRE_0(24);
ELSE
	DATA(24) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(23) <= SYNTHESIZED_WIRE_0(23);
ELSE
	DATA(23) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(22) <= SYNTHESIZED_WIRE_0(22);
ELSE
	DATA(22) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(21) <= SYNTHESIZED_WIRE_0(21);
ELSE
	DATA(21) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(20) <= SYNTHESIZED_WIRE_0(20);
ELSE
	DATA(20) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(19) <= SYNTHESIZED_WIRE_0(19);
ELSE
	DATA(19) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(18) <= SYNTHESIZED_WIRE_0(18);
ELSE
	DATA(18) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(17) <= SYNTHESIZED_WIRE_0(17);
ELSE
	DATA(17) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(16) <= SYNTHESIZED_WIRE_0(16);
ELSE
	DATA(16) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(15) <= SYNTHESIZED_WIRE_0(15);
ELSE
	DATA(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(14) <= SYNTHESIZED_WIRE_0(14);
ELSE
	DATA(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(13) <= SYNTHESIZED_WIRE_0(13);
ELSE
	DATA(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(12) <= SYNTHESIZED_WIRE_0(12);
ELSE
	DATA(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(11) <= SYNTHESIZED_WIRE_0(11);
ELSE
	DATA(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(10) <= SYNTHESIZED_WIRE_0(10);
ELSE
	DATA(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(9) <= SYNTHESIZED_WIRE_0(9);
ELSE
	DATA(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(8) <= SYNTHESIZED_WIRE_0(8);
ELSE
	DATA(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(7) <= SYNTHESIZED_WIRE_0(7);
ELSE
	DATA(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(6) <= SYNTHESIZED_WIRE_0(6);
ELSE
	DATA(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(5) <= SYNTHESIZED_WIRE_0(5);
ELSE
	DATA(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(4) <= SYNTHESIZED_WIRE_0(4);
ELSE
	DATA(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(3) <= SYNTHESIZED_WIRE_0(3);
ELSE
	DATA(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(2) <= SYNTHESIZED_WIRE_0(2);
ELSE
	DATA(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(1) <= SYNTHESIZED_WIRE_0(1);
ELSE
	DATA(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_0,SYNTHESIZED_WIRE_1)
BEGIN
if (SYNTHESIZED_WIRE_1 = '1') THEN
	DATA(0) <= SYNTHESIZED_WIRE_0(0);
ELSE
	DATA(0) <= 'Z';
END IF;
END PROCESS;


b2v_inst1 : sram32_arilla
PORT MAP(wren => wren,
		 rden => rden,
		 clock => clk,
		 address => ADDR(14 DOWNTO 2),
		 byteena => ByteEnable,
		 data => DATA,
		 q => SYNTHESIZED_WIRE_0);


HIT <= NOT(ADDR(31) OR ADDR(29) OR ADDR(30) OR ADDR(28));


PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	DFF_inst3 <= HIT;
END IF;
END PROCESS;


rden <= HIT AND RD;


wren <= HIT AND WR;


SYNTHESIZED_WIRE_1 <= DFF_inst3 AND RD;


END bdf_type;