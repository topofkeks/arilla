��l i b r a r y   i e e e ;  
 u s e   i e e e . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
 u s e   i e e e . n u m e r i c _ s t d . a l l ;  
  
 e n t i t y   S D R A M _ I n i t R O M   i s  
         p o r t (  
                 A D D R :   i n   s t d _ l o g i c _ v e c t o r ( 3   d o w n t o   0 ) ;  
                 O :   o u t   s t d _ l o g i c _ v e c t o r ( 1 1   d o w n t o   0 )  
         ) ;  
 e n d   e n t i t y ;  
  
 a r c h i t e c t u r e   r t l   o f   S D R A M _ I n i t R O M   i s  
         t y p e   r o m T y p e   i s   a r r a y   ( 1 5   d o w n t o   0 )   o f   s t d _ l o g i c _ v e c t o r ( 1 1   d o w n t o   0 ) ;  
         s i g n a l   R O M   :   r o m T y p e   : =   ( o t h e r s   = >   ( o t h e r s   = > ' 0 ' ) ) ;  
 b e g i n  
  
         - - p r o g r a m   s t a r t s   h e r e  
         R O M ( 0 ) < =   " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 1 ) < =   " 0 0 0 0 0 0 0 0 1 1 1 1 " ;  
         R O M ( 2 ) < =   " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 3 ) < =   " 0 0 0 0 0 0 0 1 0 0 1 0 " ;  
         R O M ( 4 ) < =   " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 5 ) < =   " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 6 ) < =   " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 7 ) < =   " 0 0 0 0 0 0 0 1 0 0 1 0 " ;  
         R O M ( 8 ) < =   " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 9 ) < =   " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 1 0 ) < = " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 1 1 ) < = " 0 0 0 0 0 0 1 1 0 0 1 1 " ;  
         R O M ( 1 2 ) < = " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 1 3 ) < = " 0 0 0 0 0 0 0 0 0 0 0 1 " ;  
         R O M ( 1 4 ) < = " 1 1 1 0 1 1 0 0 0 0 0 0 " ;  
         - - p r o g r a m   e n d s   h e r e  
  
 p r o c e s s ( A D D R )  
 b e g i n  
  
         O < = R O M ( t o _ i n t e g e r ( u n s i g n e d ( A D D R ) ) ) ;  
  
 e n d   p r o c e s s ;  
 e n d   r t l ;  
 