-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Sun Aug 29 03:52:12 2021"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY MemorySequencer IS 
	PORT
	(
		WR :  IN  STD_LOGIC;
		RD :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		rst :  IN  STD_LOGIC;
		color :  IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
		opX :  IN  STD_LOGIC_VECTOR(10 DOWNTO 0);
		opY :  IN  STD_LOGIC_VECTOR(10 DOWNTO 0);
		SDRAM_DQ :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		syncX :  IN  STD_LOGIC_VECTOR(10 DOWNTO 0);
		syncY :  IN  STD_LOGIC_VECTOR(10 DOWNTO 0);
		FC :  OUT  STD_LOGIC;
		O :  OUT  STD_LOGIC_VECTOR(11 DOWNTO 0);
		SDRAM_CTRL :  OUT  STD_LOGIC_VECTOR(22 DOWNTO 0)
	);
END MemorySequencer;

ARCHITECTURE bdf_type OF MemorySequencer IS 

COMPONENT mux8_14
	PORT(data0x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux8_4
	PORT(data0x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT cmp_vga_vertical
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 aeb : OUT STD_LOGIC;
		 agb : OUT STD_LOGIC;
		 alb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT const
GENERIC (const : INTEGER;
			size : INTEGER
			);
	PORT(		 data : OUT STD_LOGIC_VECTOR(size-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux2_11
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END COMPONENT;

COMPONENT cmp_vga_lastverticalline
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 aeb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cmp_vga_writeguard
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT add_vga_horizontal
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END COMPONENT;

COMPONENT cmp_vga_32readguard
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT idcreg
GENERIC (clear_value : INTEGER;
			default_value : INTEGER;
			size : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 cl : IN STD_LOGIC;
		 inc : IN STD_LOGIC;
		 dec : IN STD_LOGIC;
		 ld : IN STD_LOGIC;
		 data_in : IN STD_LOGIC_VECTOR(size-1 DOWNTO 0);
		 data_out : OUT STD_LOGIC_VECTOR(size-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT sdram_initrom
	PORT(ADDR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 O : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ldcreg
GENERIC (clear_value : INTEGER;
			default_value : INTEGER;
			size : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 cl : IN STD_LOGIC;
		 ld : IN STD_LOGIC;
		 data_in : IN STD_LOGIC_VECTOR(size-1 TO 0);
		 data_out : OUT STD_LOGIC_VECTOR(size-1 TO 0)
	);
END COMPONENT;

COMPONENT cmp_8_0
	PORT(dataa : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 aeb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cmp_vga_256readguard
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT sdram_writerom
	PORT(ADDR : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 O : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END COMPONENT;

COMPONENT cmp_vga_255
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 aeb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cmp_vga_0
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 aeb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT mux2_8
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT cmp_vga_horizontal
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 agb : OUT STD_LOGIC;
		 aleb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cmp_vga_511
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 aeb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cmp_vga_767
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 aeb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cmp_vga_799
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 aeb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT vacommandgenerator
	PORT(VA_ACT : IN STD_LOGIC;
		 VA_READ : IN STD_LOGIC;
		 VA_PRE : IN STD_LOGIC;
		 va_ADDR : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 va_Command : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dc4
	PORT(data : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 eq1 : OUT STD_LOGIC;
		 eq2 : OUT STD_LOGIC;
		 eq3 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT dc8
	PORT(data : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 eq0 : OUT STD_LOGIC;
		 eq1 : OUT STD_LOGIC;
		 eq2 : OUT STD_LOGIC;
		 eq3 : OUT STD_LOGIC;
		 eq4 : OUT STD_LOGIC;
		 eq5 : OUT STD_LOGIC;
		 eq6 : OUT STD_LOGIC;
		 eq7 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT sdram_readrom
	PORT(ADDR : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 O : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT add11
	PORT(dataa : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	actbank :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	ADDR :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	adrY :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	BA :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	CAS_N :  STD_LOGIC;
SIGNAL	CKE :  STD_LOGIC;
SIGNAL	CS_N :  STD_LOGIC;
SIGNAL	decReadCounter :  STD_LOGIC;
SIGNAL	FC_RD :  STD_LOGIC;
SIGNAL	FC_WR :  STD_LOGIC;
SIGNAL	first_read :  STD_LOGIC;
SIGNAL	FREE_RANGE :  STD_LOGIC;
SIGNAL	HORIZONTAL_FREE_RANGE :  STD_LOGIC;
SIGNAL	HORIZONTAL_VISIBLE_AREA :  STD_LOGIC;
SIGNAL	init_ADDR :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	init_Command :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	initrom_ba :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	initrom_bruncnd :  STD_LOGIC;
SIGNAL	last_line :  STD_LOGIC;
SIGNAL	lastBank :  STD_LOGIC;
SIGNAL	ldReadCounter :  STD_LOGIC;
SIGNAL	memX :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	memY :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	no_read :  STD_LOGIC;
SIGNAL	no_write :  STD_LOGIC;
SIGNAL	one :  STD_LOGIC;
SIGNAL	pre_bank :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	RAS_N :  STD_LOGIC;
SIGNAL	rd256_guard :  STD_LOGIC;
SIGNAL	rd32_guard :  STD_LOGIC;
SIGNAL	rd_ADDR :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	RD_BUS :  STD_LOGIC;
SIGNAL	rd_Command :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	RDreq :  STD_LOGIC;
SIGNAL	read_guard :  STD_LOGIC;
SIGNAL	readComplete :  STD_LOGIC;
SIGNAL	readrom_ba :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	readrom_cc :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	ready :  STD_LOGIC;
SIGNAL	va_ADDR :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	va_Command :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	VERTICAL_FREE_RANGE :  STD_LOGIC;
SIGNAL	VERTICAL_VISIBLE_AREA :  STD_LOGIC;
SIGNAL	VERTICAL_VISIBLE_EXCEPT_LAST :  STD_LOGIC;
SIGNAL	VISIBLE_AREA :  STD_LOGIC;
SIGNAL	WE_N :  STD_LOGIC;
SIGNAL	wr_ADDR :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	WR_BUS :  STD_LOGIC;
SIGNAL	wr_Command :  STD_LOGIC_VECTOR(2 DOWNTO 1);
SIGNAL	write_guard :  STD_LOGIC;
SIGNAL	writerom_ba :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	writerom_brno_write :  STD_LOGIC;
SIGNAL	writerom_brnot_ready :  STD_LOGIC;
SIGNAL	writerom_bruncnd :  STD_LOGIC;
SIGNAL	writerom_cc :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	WRreq :  STD_LOGIC;
SIGNAL	zero :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC_VECTOR(10 DOWNTO 0);

SIGNAL	GDFX_TEMP_SIGNAL_25 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_20 :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_18 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_17 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_8 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_19 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_6 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_5 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_7 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_23 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_27 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_22 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_28 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_24 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_26 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_21 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_29 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_14 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_16 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_15 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_13 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_12 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_11 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_10 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_9 :  STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN 

readrom_ba(2) <= GDFX_TEMP_SIGNAL_25(15);
readrom_ba(1) <= GDFX_TEMP_SIGNAL_25(14);
readrom_ba(0) <= GDFX_TEMP_SIGNAL_25(13);
readrom_cc(2) <= GDFX_TEMP_SIGNAL_25(12);
readrom_cc(1) <= GDFX_TEMP_SIGNAL_25(11);
readrom_cc(0) <= GDFX_TEMP_SIGNAL_25(10);
rd_Command(2) <= GDFX_TEMP_SIGNAL_25(9);
decReadCounter <= GDFX_TEMP_SIGNAL_25(8);
RD_BUS <= GDFX_TEMP_SIGNAL_25(7);
FC_RD <= GDFX_TEMP_SIGNAL_25(6);
ldReadCounter <= GDFX_TEMP_SIGNAL_25(5);
rd_ADDR(1) <= GDFX_TEMP_SIGNAL_25(4);
rd_Command(0) <= GDFX_TEMP_SIGNAL_25(3);
rd_ADDR(0) <= GDFX_TEMP_SIGNAL_25(2);
rd_ADDR(2) <= GDFX_TEMP_SIGNAL_25(1);
rd_Command(1) <= GDFX_TEMP_SIGNAL_25(0);

writerom_ba(2) <= GDFX_TEMP_SIGNAL_20(10);
writerom_ba(1) <= GDFX_TEMP_SIGNAL_20(9);
writerom_ba(0) <= GDFX_TEMP_SIGNAL_20(8);
writerom_cc(1) <= GDFX_TEMP_SIGNAL_20(7);
writerom_cc(0) <= GDFX_TEMP_SIGNAL_20(6);
WR_BUS <= GDFX_TEMP_SIGNAL_20(5);
wr_ADDR(1) <= GDFX_TEMP_SIGNAL_20(4);
wr_Command(2) <= GDFX_TEMP_SIGNAL_20(3);
wr_ADDR(2) <= GDFX_TEMP_SIGNAL_20(2);
wr_Command(1) <= GDFX_TEMP_SIGNAL_20(1);

initrom_ba(3) <= GDFX_TEMP_SIGNAL_18(11);
initrom_ba(2) <= GDFX_TEMP_SIGNAL_18(10);
initrom_ba(1) <= GDFX_TEMP_SIGNAL_18(9);
initrom_ba(0) <= GDFX_TEMP_SIGNAL_18(8);
initrom_bruncnd <= GDFX_TEMP_SIGNAL_18(7);
ready <= GDFX_TEMP_SIGNAL_18(6);
init_ADDR(2) <= GDFX_TEMP_SIGNAL_18(5);
init_Command(1) <= GDFX_TEMP_SIGNAL_18(4);
init_ADDR(0) <= GDFX_TEMP_SIGNAL_18(3);
init_ADDR(1) <= GDFX_TEMP_SIGNAL_18(2);
init_Command(2) <= GDFX_TEMP_SIGNAL_18(1);
init_Command(0) <= GDFX_TEMP_SIGNAL_18(0);

CS_N <= GDFX_TEMP_SIGNAL_17(3);
RAS_N <= GDFX_TEMP_SIGNAL_17(2);
CAS_N <= GDFX_TEMP_SIGNAL_17(1);
WE_N <= GDFX_TEMP_SIGNAL_17(0);

BA(1) <= GDFX_TEMP_SIGNAL_8(13);
BA(0) <= GDFX_TEMP_SIGNAL_8(12);
ADDR(11) <= GDFX_TEMP_SIGNAL_8(11);
ADDR(10) <= GDFX_TEMP_SIGNAL_8(10);
ADDR(9) <= GDFX_TEMP_SIGNAL_8(9);
ADDR(8) <= GDFX_TEMP_SIGNAL_8(8);
ADDR(7) <= GDFX_TEMP_SIGNAL_8(7);
ADDR(6) <= GDFX_TEMP_SIGNAL_8(6);
ADDR(5) <= GDFX_TEMP_SIGNAL_8(5);
ADDR(4) <= GDFX_TEMP_SIGNAL_8(4);
ADDR(3) <= GDFX_TEMP_SIGNAL_8(3);
ADDR(2) <= GDFX_TEMP_SIGNAL_8(2);
ADDR(1) <= GDFX_TEMP_SIGNAL_8(1);
ADDR(0) <= GDFX_TEMP_SIGNAL_8(0);

GDFX_TEMP_SIGNAL_1 <= (actbank(1 DOWNTO 0) & zero & adrY(10 DOWNTO 0));
GDFX_TEMP_SIGNAL_2 <= (actbank(1 DOWNTO 0) & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero);
GDFX_TEMP_SIGNAL_19 <= (wr_Command(2 DOWNTO 1) & zero);
GDFX_TEMP_SIGNAL_3 <= (opX(9 DOWNTO 8) & zero & one & zero & zero & opX(7 DOWNTO 0));
GDFX_TEMP_SIGNAL_6 <= (opX(9 DOWNTO 8) & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero);
GDFX_TEMP_SIGNAL_5 <= (opX(9 DOWNTO 8) & zero & opY(10 DOWNTO 0));
GDFX_TEMP_SIGNAL_7 <= (pre_bank(1 DOWNTO 0) & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero);
GDFX_TEMP_SIGNAL_4 <= (zero & zero & zero & zero & one & zero & zero & zero & one & zero & zero & one & one & one);
GDFX_TEMP_SIGNAL_0 <= (zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero & zero);
GDFX_TEMP_SIGNAL_23 <= (one & zero);
GDFX_TEMP_SIGNAL_27 <= (one & zero);
GDFX_TEMP_SIGNAL_22 <= (zero & one);
GDFX_TEMP_SIGNAL_28 <= (zero & one);
GDFX_TEMP_SIGNAL_24 <= (one & one);
GDFX_TEMP_SIGNAL_26 <= (one & one);
GDFX_TEMP_SIGNAL_21 <= (zero & zero);
GDFX_TEMP_SIGNAL_29 <= (zero & zero);
GDFX_TEMP_SIGNAL_14 <= (zero & zero & one & zero);
GDFX_TEMP_SIGNAL_16 <= (zero & zero & zero & zero);
GDFX_TEMP_SIGNAL_15 <= (zero & zero & zero & one);
GDFX_TEMP_SIGNAL_13 <= (zero & one & zero & zero);
GDFX_TEMP_SIGNAL_12 <= (zero & one & zero & one);
GDFX_TEMP_SIGNAL_11 <= (zero & zero & one & one);
GDFX_TEMP_SIGNAL_10 <= (zero & one & one & one);
GDFX_TEMP_SIGNAL_9 <= (one & zero & zero & zero);


b2v_AddressMux : mux8_14
PORT MAP(data0x => GDFX_TEMP_SIGNAL_0,
		 data1x => GDFX_TEMP_SIGNAL_1,
		 data2x => GDFX_TEMP_SIGNAL_2,
		 data3x => GDFX_TEMP_SIGNAL_3,
		 data4x => GDFX_TEMP_SIGNAL_4,
		 data5x => GDFX_TEMP_SIGNAL_5,
		 data6x => GDFX_TEMP_SIGNAL_6,
		 data7x => GDFX_TEMP_SIGNAL_7,
		 sel => SYNTHESIZED_WIRE_0,
		 result => GDFX_TEMP_SIGNAL_8);


b2v_CommandMux : mux8_4
PORT MAP(data0x => GDFX_TEMP_SIGNAL_9,
		 data1x => GDFX_TEMP_SIGNAL_10,
		 data2x => GDFX_TEMP_SIGNAL_11,
		 data3x => GDFX_TEMP_SIGNAL_12,
		 data4x => GDFX_TEMP_SIGNAL_13,
		 data5x => GDFX_TEMP_SIGNAL_14,
		 data6x => GDFX_TEMP_SIGNAL_15,
		 data7x => GDFX_TEMP_SIGNAL_16,
		 sel => SYNTHESIZED_WIRE_1,
		 result => GDFX_TEMP_SIGNAL_17);


b2v_inst : cmp_vga_vertical
PORT MAP(dataa => memY,
		 aeb => SYNTHESIZED_WIRE_64,
		 alb => VERTICAL_VISIBLE_EXCEPT_LAST);

memY <= syncY;




b2v_inst100 : const
GENERIC MAP(const => 1,
			size => 11
			)
PORT MAP(		 data => SYNTHESIZED_WIRE_65);


SYNTHESIZED_WIRE_51 <= HORIZONTAL_VISIBLE_AREA AND VERTICAL_VISIBLE_AREA;


b2v_inst102 : mux2_11
PORT MAP(sel => last_line,
		 data0x => SYNTHESIZED_WIRE_2,
		 data1x => SYNTHESIZED_WIRE_3,
		 result => adrY);


b2v_inst103 : const
GENERIC MAP(const => 0,
			size => 11
			)
PORT MAP(		 data => SYNTHESIZED_WIRE_3);



b2v_inst12 : cmp_vga_lastverticalline
PORT MAP(dataa => memY,
		 aeb => last_line);


b2v_inst13 : cmp_vga_writeguard
PORT MAP(dataa => memX,
		 ageb => write_guard);


b2v_inst14 : add_vga_horizontal
PORT MAP(dataa => syncX,
		 result => memX);


SYNTHESIZED_WIRE_0 <= init_ADDR OR wr_ADDR OR rd_ADDR OR va_ADDR;

CKE <= one;



b2v_inst17 : cmp_vga_32readguard
PORT MAP(dataa => memX,
		 ageb => rd32_guard);


b2v_inst18 : idcreg
GENERIC MAP(clear_value => 0,
			default_value => 0,
			size => 4
			)
PORT MAP(clk => clk,
		 cl => rst,
		 inc => one,
		 dec => zero,
		 ld => initrom_bruncnd,
		 data_in => initrom_ba,
		 data_out => SYNTHESIZED_WIRE_4);


b2v_inst19 : sdram_initrom
PORT MAP(ADDR => SYNTHESIZED_WIRE_4,
		 O => GDFX_TEMP_SIGNAL_18);


b2v_inst2 : ldcreg
GENERIC MAP(clear_value => 0,
			default_value => 0,
			size => 1
			)
PORT MAP(clk => clk,
		 cl => WR_BUS,
		 ld => WR,
		 data_in(0) => one,
		 data_out(0) => WRreq);


SYNTHESIZED_WIRE_1 <= init_Command OR GDFX_TEMP_SIGNAL_19 OR rd_Command OR va_Command;


b2v_inst21 : cmp_8_0
PORT MAP(dataa => SYNTHESIZED_WIRE_5,
		 aeb => readComplete);


b2v_inst22 : cmp_vga_256readguard
PORT MAP(dataa => memX,
		 ageb => rd256_guard);


b2v_inst23 : sdram_writerom
PORT MAP(ADDR => SYNTHESIZED_WIRE_6,
		 O => GDFX_TEMP_SIGNAL_20);


b2v_inst24 : cmp_vga_255
PORT MAP(dataa => memX,
		 aeb => SYNTHESIZED_WIRE_32);


b2v_inst25 : cmp_vga_0
PORT MAP(dataa => memX,
		 aeb => first_read);


b2v_inst26 : mux2_8
PORT MAP(sel => lastBank,
		 data0x => SYNTHESIZED_WIRE_7,
		 data1x => SYNTHESIZED_WIRE_8,
		 result => SYNTHESIZED_WIRE_58);


lastBank <= opX(9) AND opX(8);


b2v_inst28 : const
GENERIC MAP(const => 30,
			size => 8
			)
PORT MAP(		 data => SYNTHESIZED_WIRE_8);


SYNTHESIZED_WIRE_78 <= SYNTHESIZED_WIRE_9 AND VISIBLE_AREA;


b2v_inst3 : cmp_vga_horizontal
PORT MAP(dataa => memX,
		 aleb => HORIZONTAL_VISIBLE_AREA);


SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_10 AND VISIBLE_AREA;


SYNTHESIZED_WIRE_68 <= SYNTHESIZED_WIRE_11 AND VISIBLE_AREA;


b2v_inst33 : cmp_vga_511
PORT MAP(dataa => memX,
		 aeb => SYNTHESIZED_WIRE_11);


b2v_inst34 : cmp_vga_767
PORT MAP(dataa => memX,
		 aeb => SYNTHESIZED_WIRE_10);


b2v_inst35 : cmp_vga_799
PORT MAP(dataa => memX,
		 aeb => SYNTHESIZED_WIRE_9);


b2v_inst36 : vacommandgenerator
PORT MAP(VA_ACT => SYNTHESIZED_WIRE_12,
		 VA_READ => SYNTHESIZED_WIRE_13,
		 VA_PRE => SYNTHESIZED_WIRE_14,
		 va_ADDR => va_ADDR,
		 va_Command => va_Command);


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_67 OR SYNTHESIZED_WIRE_68 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_70;


b2v_inst38 : idcreg
GENERIC MAP(clear_value => 0,
			default_value => 0,
			size => 3
			)
PORT MAP(clk => clk,
		 cl => rst,
		 inc => one,
		 dec => zero,
		 ld => SYNTHESIZED_WIRE_19,
		 data_in => writerom_ba,
		 data_out => SYNTHESIZED_WIRE_6);


b2v_inst39 : dc4
PORT MAP(data => writerom_cc,
		 eq1 => writerom_bruncnd,
		 eq2 => writerom_brnot_ready,
		 eq3 => writerom_brno_write);


wr_ADDR(0) <= wr_ADDR(1) OR wr_ADDR(2);


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_20 OR SYNTHESIZED_WIRE_21 OR writerom_bruncnd;


SYNTHESIZED_WIRE_20 <= writerom_brnot_ready AND SYNTHESIZED_WIRE_22;


SYNTHESIZED_WIRE_21 <= writerom_brno_write AND no_write;


SYNTHESIZED_WIRE_75 <= VERTICAL_VISIBLE_AREA AND HORIZONTAL_VISIBLE_AREA;


SYNTHESIZED_WIRE_26 <= VERTICAL_VISIBLE_AREA AND write_guard;


SYNTHESIZED_WIRE_24 <= last_line AND write_guard;


SYNTHESIZED_WIRE_22 <= NOT(ready);



SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_71 OR SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_73 OR SYNTHESIZED_WIRE_74;


no_write <= SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_24 OR SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_25 <= NOT(WRreq);

O<= syncY(1 downto 0) & syncX(9 downto 0);


PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(11) <= color(11);
ELSE
	SDRAM_DQ(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(10) <= color(10);
ELSE
	SDRAM_DQ(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(9) <= color(9);
ELSE
	SDRAM_DQ(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(8) <= color(8);
ELSE
	SDRAM_DQ(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(7) <= color(7);
ELSE
	SDRAM_DQ(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(6) <= color(6);
ELSE
	SDRAM_DQ(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(5) <= color(5);
ELSE
	SDRAM_DQ(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(4) <= color(4);
ELSE
	SDRAM_DQ(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(3) <= color(3);
ELSE
	SDRAM_DQ(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(2) <= color(2);
ELSE
	SDRAM_DQ(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(1) <= color(1);
ELSE
	SDRAM_DQ(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(color,WR_BUS)
BEGIN
if (WR_BUS = '1') THEN
	SDRAM_DQ(0) <= color(0);
ELSE
	SDRAM_DQ(0) <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_14 <= SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_77 OR SYNTHESIZED_WIRE_78 OR SYNTHESIZED_WIRE_79;


b2v_inst53 : const
GENERIC MAP(const => 254,
			size => 8
			)
PORT MAP(		 data => SYNTHESIZED_WIRE_7);


no_read <= zero OR SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29 OR WRreq OR SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_75;


SYNTHESIZED_WIRE_70 <= SYNTHESIZED_WIRE_32 AND VISIBLE_AREA;


SYNTHESIZED_WIRE_67 <= first_read AND SYNTHESIZED_WIRE_33;


PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_71 <= SYNTHESIZED_WIRE_67;
END IF;
END PROCESS;


PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_74 <= SYNTHESIZED_WIRE_70;
END IF;
END PROCESS;


PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_76 <= SYNTHESIZED_WIRE_74;
END IF;
END PROCESS;



PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_72 <= SYNTHESIZED_WIRE_68;
END IF;
END PROCESS;


PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_79 <= SYNTHESIZED_WIRE_72;
END IF;
END PROCESS;


PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_69;
END IF;
END PROCESS;


PROCESS(clk)
BEGIN
IF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_77 <= SYNTHESIZED_WIRE_73;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_30 <= NOT(RDreq);



PROCESS(GDFX_TEMP_SIGNAL_21,SYNTHESIZED_WIRE_76)
BEGIN
if (SYNTHESIZED_WIRE_76 = '1') THEN
	pre_bank(1) <= GDFX_TEMP_SIGNAL_21(1);
ELSE
	pre_bank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_21,SYNTHESIZED_WIRE_76)
BEGIN
if (SYNTHESIZED_WIRE_76 = '1') THEN
	pre_bank(0) <= GDFX_TEMP_SIGNAL_21(0);
ELSE
	pre_bank(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(GDFX_TEMP_SIGNAL_22,SYNTHESIZED_WIRE_79)
BEGIN
if (SYNTHESIZED_WIRE_79 = '1') THEN
	pre_bank(1) <= GDFX_TEMP_SIGNAL_22(1);
ELSE
	pre_bank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_22,SYNTHESIZED_WIRE_79)
BEGIN
if (SYNTHESIZED_WIRE_79 = '1') THEN
	pre_bank(0) <= GDFX_TEMP_SIGNAL_22(0);
ELSE
	pre_bank(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(GDFX_TEMP_SIGNAL_23,SYNTHESIZED_WIRE_77)
BEGIN
if (SYNTHESIZED_WIRE_77 = '1') THEN
	pre_bank(1) <= GDFX_TEMP_SIGNAL_23(1);
ELSE
	pre_bank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_23,SYNTHESIZED_WIRE_77)
BEGIN
if (SYNTHESIZED_WIRE_77 = '1') THEN
	pre_bank(0) <= GDFX_TEMP_SIGNAL_23(0);
ELSE
	pre_bank(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(GDFX_TEMP_SIGNAL_24,SYNTHESIZED_WIRE_78)
BEGIN
if (SYNTHESIZED_WIRE_78 = '1') THEN
	pre_bank(1) <= GDFX_TEMP_SIGNAL_24(1);
ELSE
	pre_bank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_24,SYNTHESIZED_WIRE_78)
BEGIN
if (SYNTHESIZED_WIRE_78 = '1') THEN
	pre_bank(0) <= GDFX_TEMP_SIGNAL_24(0);
ELSE
	pre_bank(0) <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_42 <= rd32_guard AND lastBank;


SYNTHESIZED_WIRE_41 <= rd256_guard AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_40 <= NOT(lastBank);



read_guard <= SYNTHESIZED_WIRE_41 OR SYNTHESIZED_WIRE_42;


SYNTHESIZED_WIRE_28 <= read_guard AND last_line;


SYNTHESIZED_WIRE_29 <= VERTICAL_VISIBLE_AREA AND read_guard;


b2v_inst75 : dc8
PORT MAP(data => readrom_cc,
		 eq1 => SYNTHESIZED_WIRE_47,
		 eq2 => SYNTHESIZED_WIRE_49,
		 eq3 => SYNTHESIZED_WIRE_52,
		 eq4 => SYNTHESIZED_WIRE_53);


b2v_inst76 : idcreg
GENERIC MAP(clear_value => 0,
			default_value => 0,
			size => 3
			)
PORT MAP(clk => clk,
		 cl => rst,
		 inc => one,
		 dec => zero,
		 ld => SYNTHESIZED_WIRE_43,
		 data_in => readrom_ba,
		 data_out => SYNTHESIZED_WIRE_44);


b2v_inst77 : sdram_readrom
PORT MAP(ADDR => SYNTHESIZED_WIRE_44,
		 O => GDFX_TEMP_SIGNAL_25);


SYNTHESIZED_WIRE_43 <= SYNTHESIZED_WIRE_45 OR SYNTHESIZED_WIRE_46 OR SYNTHESIZED_WIRE_47 OR SYNTHESIZED_WIRE_48;


SYNTHESIZED_WIRE_45 <= SYNTHESIZED_WIRE_49 AND SYNTHESIZED_WIRE_50;


VISIBLE_AREA <= SYNTHESIZED_WIRE_51 AND ready;


SYNTHESIZED_WIRE_50 <= NOT(ready);



SYNTHESIZED_WIRE_48 <= SYNTHESIZED_WIRE_52 AND no_read;


SYNTHESIZED_WIRE_46 <= SYNTHESIZED_WIRE_53 AND SYNTHESIZED_WIRE_54;


SYNTHESIZED_WIRE_54 <= NOT(readComplete);



FC <= FC_RD OR WR_BUS;

RDreq <= RD;



PROCESS(GDFX_TEMP_SIGNAL_26,SYNTHESIZED_WIRE_55)
BEGIN
if (SYNTHESIZED_WIRE_55 = '1') THEN
	actbank(1) <= GDFX_TEMP_SIGNAL_26(1);
ELSE
	actbank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_26,SYNTHESIZED_WIRE_55)
BEGIN
if (SYNTHESIZED_WIRE_55 = '1') THEN
	actbank(0) <= GDFX_TEMP_SIGNAL_26(0);
ELSE
	actbank(0) <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_33 <= VERTICAL_VISIBLE_EXCEPT_LAST OR last_line;


PROCESS(GDFX_TEMP_SIGNAL_27,SYNTHESIZED_WIRE_56)
BEGIN
if (SYNTHESIZED_WIRE_56 = '1') THEN
	actbank(1) <= GDFX_TEMP_SIGNAL_27(1);
ELSE
	actbank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_27,SYNTHESIZED_WIRE_56)
BEGIN
if (SYNTHESIZED_WIRE_56 = '1') THEN
	actbank(0) <= GDFX_TEMP_SIGNAL_27(0);
ELSE
	actbank(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(GDFX_TEMP_SIGNAL_28,SYNTHESIZED_WIRE_57)
BEGIN
if (SYNTHESIZED_WIRE_57 = '1') THEN
	actbank(1) <= GDFX_TEMP_SIGNAL_28(1);
ELSE
	actbank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_28,SYNTHESIZED_WIRE_57)
BEGIN
if (SYNTHESIZED_WIRE_57 = '1') THEN
	actbank(0) <= GDFX_TEMP_SIGNAL_28(0);
ELSE
	actbank(0) <= 'Z';
END IF;
END PROCESS;


b2v_inst9 : idcreg
GENERIC MAP(clear_value => 0,
			default_value => 0,
			size => 8
			)
PORT MAP(clk => clk,
		 cl => zero,
		 inc => zero,
		 dec => decReadCounter,
		 ld => ldReadCounter,
		 data_in => SYNTHESIZED_WIRE_58,
		 data_out => SYNTHESIZED_WIRE_5);


PROCESS(GDFX_TEMP_SIGNAL_29,SYNTHESIZED_WIRE_59)
BEGIN
if (SYNTHESIZED_WIRE_59 = '1') THEN
	actbank(1) <= GDFX_TEMP_SIGNAL_29(1);
ELSE
	actbank(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(GDFX_TEMP_SIGNAL_29,SYNTHESIZED_WIRE_59)
BEGIN
if (SYNTHESIZED_WIRE_59 = '1') THEN
	actbank(0) <= GDFX_TEMP_SIGNAL_29(0);
ELSE
	actbank(0) <= 'Z';
END IF;
END PROCESS;


SYNTHESIZED_WIRE_55 <= SYNTHESIZED_WIRE_73 OR SYNTHESIZED_WIRE_69;


SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_59 <= SYNTHESIZED_WIRE_71 OR SYNTHESIZED_WIRE_67;


SYNTHESIZED_WIRE_57 <= SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_70;


VERTICAL_VISIBLE_AREA <= VERTICAL_VISIBLE_EXCEPT_LAST OR SYNTHESIZED_WIRE_64;


b2v_inst98 : add11
PORT MAP(dataa => SYNTHESIZED_WIRE_65,
		 datab => memY,
		 result => SYNTHESIZED_WIRE_66);


b2v_inst99 : mux2_11
PORT MAP(sel => first_read,
		 data0x => memY,
		 data1x => SYNTHESIZED_WIRE_66,
		 result => SYNTHESIZED_WIRE_2);

SDRAM_CTRL(22) <= zero;
SDRAM_CTRL(21 DOWNTO 10) <= ADDR;
SDRAM_CTRL(9 DOWNTO 8) <= BA;
SDRAM_CTRL(7) <= RAS_N;
SDRAM_CTRL(6) <= CAS_N;
SDRAM_CTRL(5) <= zero;
SDRAM_CTRL(4) <= zero;
SDRAM_CTRL(3) <= CKE;
SDRAM_CTRL(2) <= clk;
SDRAM_CTRL(1) <= WE_N;
SDRAM_CTRL(0) <= CS_N;

ADDR(11 DOWNTO 0) <= GDFX_TEMP_SIGNAL_8(11 DOWNTO 0);
BA(1 DOWNTO 0) <= GDFX_TEMP_SIGNAL_8(13 DOWNTO 12);
CAS_N <= GDFX_TEMP_SIGNAL_17(1);
CS_N <= GDFX_TEMP_SIGNAL_17(3);
decReadCounter <= GDFX_TEMP_SIGNAL_25(8);
FC_RD <= GDFX_TEMP_SIGNAL_25(6);
FC_WR <= GDFX_TEMP_SIGNAL_20(2);
initrom_ba(3 DOWNTO 0) <= GDFX_TEMP_SIGNAL_18(11 DOWNTO 8);
initrom_bruncnd <= GDFX_TEMP_SIGNAL_18(7);
ldReadCounter <= GDFX_TEMP_SIGNAL_25(5);
one <= '1';
RAS_N <= GDFX_TEMP_SIGNAL_17(2);
RD_BUS <= GDFX_TEMP_SIGNAL_25(7);
readrom_ba(2 DOWNTO 0) <= GDFX_TEMP_SIGNAL_25(15 DOWNTO 13);
readrom_cc(2 DOWNTO 0) <= GDFX_TEMP_SIGNAL_25(12 DOWNTO 10);
ready <= GDFX_TEMP_SIGNAL_18(6);
WE_N <= GDFX_TEMP_SIGNAL_17(0);
WR_BUS <= GDFX_TEMP_SIGNAL_20(5);
writerom_ba(2 DOWNTO 0) <= GDFX_TEMP_SIGNAL_20(10 DOWNTO 8);
writerom_cc(1 DOWNTO 0) <= GDFX_TEMP_SIGNAL_20(7 DOWNTO 6);
zero <= '0';
END bdf_type;